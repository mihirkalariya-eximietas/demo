sfaf
sdgsdg
