sdjbsi
adgs
